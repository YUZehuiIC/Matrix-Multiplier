
module MatrixMultiplier ( CLK, NRST, START, A, B, OUT, OUT_STROBE );
  input [7:0] A;
  input [7:0] B;
  output [16:0] OUT;
  input CLK, NRST, START;
  output OUT_STROBE;
  wire   \next_state[1] , N13, N14, N15, N16, N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, P_temp_16, \P_temp[9] , \P_temp[8] , \P_temp[7] , \P_temp[6] ,
         \P_temp[5] , \P_temp[4] , \P_temp[3] , \P_temp[2] , \P_temp[1] ,
         \P_temp[14] , \P_temp[13] , \P_temp[12] , \P_temp[11] , \P_temp[10] ,
         \P_temp[0] , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159;
  wire   [1:0] state;
  wire   [16:0] Add2;

  TFEP3 Flag_reg ( .T(n60), .C(CLK), .SN(n154), .QN(n19) );
  DFC3 \Add2_reg[16]  ( .D(n131), .C(CLK), .RN(NRST), .Q(Add2[16]), .QN(n2) );
  DFC3 \Add2_reg[15]  ( .D(n129), .C(CLK), .RN(NRST), .Q(Add2[15]), .QN(n3) );
  DFC3 \Add2_reg[14]  ( .D(n127), .C(CLK), .RN(NRST), .Q(Add2[14]), .QN(n4) );
  DFC3 \Add2_reg[13]  ( .D(n125), .C(CLK), .RN(NRST), .Q(Add2[13]), .QN(n5) );
  DFC3 \Add2_reg[12]  ( .D(n123), .C(CLK), .RN(NRST), .Q(Add2[12]), .QN(n6) );
  DFC3 \Add2_reg[11]  ( .D(n121), .C(CLK), .RN(NRST), .Q(Add2[11]), .QN(n7) );
  DFC3 \Add2_reg[10]  ( .D(n119), .C(CLK), .RN(NRST), .Q(Add2[10]), .QN(n8) );
  DFC3 \Add2_reg[9]  ( .D(n117), .C(CLK), .RN(NRST), .Q(Add2[9]), .QN(n9) );
  DFC3 \Add2_reg[8]  ( .D(n115), .C(CLK), .RN(NRST), .Q(Add2[8]), .QN(n10) );
  DFC3 \Add2_reg[7]  ( .D(n113), .C(CLK), .RN(NRST), .Q(Add2[7]), .QN(n11) );
  DFC3 \Add2_reg[6]  ( .D(n111), .C(CLK), .RN(NRST), .Q(Add2[6]), .QN(n12) );
  DFC3 \Add2_reg[5]  ( .D(n109), .C(CLK), .RN(NRST), .Q(Add2[5]), .QN(n13) );
  DFC3 \Add2_reg[4]  ( .D(n107), .C(CLK), .RN(NRST), .Q(Add2[4]), .QN(n14) );
  DFC3 \Add2_reg[3]  ( .D(n105), .C(CLK), .RN(NRST), .Q(Add2[3]), .QN(n15) );
  DFC3 \Add2_reg[2]  ( .D(n103), .C(CLK), .RN(NRST), .Q(Add2[2]), .QN(n16) );
  DFC3 \Add2_reg[1]  ( .D(n101), .C(CLK), .RN(NRST), .Q(Add2[1]), .QN(n17) );
  DFC3 \Add2_reg[0]  ( .D(n99), .C(CLK), .RN(NRST), .Q(Add2[0]), .QN(n18) );
  OAI212 U4 ( .A(n42), .B(n20), .C(n43), .Q(n64) );
  OAI212 U6 ( .A(n42), .B(n21), .C(n44), .Q(n65) );
  OAI212 U8 ( .A(n42), .B(n22), .C(n45), .Q(n66) );
  OAI212 U10 ( .A(n153), .B(n23), .C(n46), .Q(n67) );
  OAI212 U12 ( .A(n42), .B(n24), .C(n47), .Q(n68) );
  OAI212 U14 ( .A(n42), .B(n25), .C(n48), .Q(n69) );
  OAI212 U16 ( .A(n42), .B(n26), .C(n49), .Q(n70) );
  OAI212 U18 ( .A(n42), .B(n27), .C(n50), .Q(n71) );
  OAI212 U20 ( .A(n42), .B(n28), .C(n51), .Q(n72) );
  OAI212 U22 ( .A(n42), .B(n29), .C(n52), .Q(n73) );
  OAI212 U24 ( .A(n42), .B(n30), .C(n53), .Q(n74) );
  OAI212 U26 ( .A(n42), .B(n31), .C(n54), .Q(n75) );
  OAI212 U28 ( .A(n153), .B(n32), .C(n55), .Q(n76) );
  OAI212 U30 ( .A(n153), .B(n33), .C(n56), .Q(n77) );
  OAI212 U32 ( .A(n153), .B(n34), .C(n57), .Q(n78) );
  OAI212 U34 ( .A(n153), .B(n35), .C(n58), .Q(n79) );
  OAI212 U36 ( .A(n153), .B(n36), .C(n59), .Q(n80) );
  DFC3 \state_reg[0]  ( .D(n156), .C(CLK), .RN(NRST), .Q(state[0]), .QN(n40)
         );
  TFEC3 \state_reg[1]  ( .T(n152), .C(CLK), .RN(NRST), .Q(state[1]) );
  DFC3 \OUT_reg[16]  ( .D(n151), .C(CLK), .RN(n154), .Q(OUT[16]) );
  DFC3 \OUT_reg[15]  ( .D(n150), .C(CLK), .RN(n154), .Q(OUT[15]) );
  DFC3 \OUT_reg[14]  ( .D(n149), .C(CLK), .RN(n154), .Q(OUT[14]) );
  DFC3 \OUT_reg[13]  ( .D(n148), .C(CLK), .RN(n154), .Q(OUT[13]) );
  DFC3 \OUT_reg[12]  ( .D(n147), .C(CLK), .RN(n154), .Q(OUT[12]) );
  DFC3 \OUT_reg[11]  ( .D(n146), .C(CLK), .RN(n154), .Q(OUT[11]) );
  DFC3 \OUT_reg[10]  ( .D(n145), .C(CLK), .RN(n154), .Q(OUT[10]) );
  DFC3 \OUT_reg[9]  ( .D(n144), .C(CLK), .RN(n154), .Q(OUT[9]) );
  DFC3 \OUT_reg[8]  ( .D(n143), .C(CLK), .RN(n154), .Q(OUT[8]) );
  DFC3 \OUT_reg[7]  ( .D(n142), .C(CLK), .RN(NRST), .Q(OUT[7]) );
  DFC3 \OUT_reg[6]  ( .D(n141), .C(CLK), .RN(n155), .Q(OUT[6]) );
  DFC3 \OUT_reg[5]  ( .D(n140), .C(CLK), .RN(NRST), .Q(OUT[5]) );
  DFC3 \OUT_reg[4]  ( .D(n139), .C(CLK), .RN(n154), .Q(OUT[4]) );
  DFC3 \OUT_reg[3]  ( .D(n138), .C(CLK), .RN(n155), .Q(OUT[3]) );
  DFC3 \OUT_reg[2]  ( .D(n137), .C(CLK), .RN(n154), .Q(OUT[2]) );
  DFC3 \OUT_reg[1]  ( .D(n136), .C(CLK), .RN(n155), .Q(OUT[1]) );
  DFC3 \OUT_reg[0]  ( .D(n135), .C(CLK), .RN(NRST), .Q(OUT[0]) );
  MatrixMultiplier_DW_mult_tc_0 mult_38 ( .a(A), .b(B), .product({P_temp_16, 
        \P_temp[14] , \P_temp[13] , \P_temp[12] , \P_temp[11] , \P_temp[10] , 
        \P_temp[9] , \P_temp[8] , \P_temp[7] , \P_temp[6] , \P_temp[5] , 
        \P_temp[4] , \P_temp[3] , \P_temp[2] , \P_temp[1] , \P_temp[0] }) );
  MatrixMultiplier_DW01_add_0 add_53 ( .A({P_temp_16, P_temp_16, \P_temp[14] , 
        \P_temp[13] , \P_temp[12] , \P_temp[11] , \P_temp[10] , \P_temp[9] , 
        \P_temp[8] , \P_temp[7] , \P_temp[6] , \P_temp[5] , \P_temp[4] , 
        \P_temp[3] , \P_temp[2] , \P_temp[1] , \P_temp[0] }), .B({Add2[16:1], 
        n134}), .CI(n159), .SUM({N29, N28, N27, N26, N25, N24, N23, N22, N21, 
        N20, N19, N18, N17, N16, N15, N14, N13}) );
  DFEC1 \Addsum_reg[16]  ( .D(N29), .E(n63), .C(CLK), .RN(NRST), .QN(n20) );
  DFEC1 \Addsum_reg[15]  ( .D(N28), .E(n63), .C(CLK), .RN(NRST), .QN(n21) );
  DFEC1 \Addsum_reg[14]  ( .D(N27), .E(n63), .C(CLK), .RN(NRST), .QN(n22) );
  DFEC1 \Addsum_reg[13]  ( .D(N26), .E(n63), .C(CLK), .RN(NRST), .QN(n23) );
  DFEC1 \Addsum_reg[12]  ( .D(N25), .E(n63), .C(CLK), .RN(NRST), .QN(n24) );
  DFEC1 \Addsum_reg[11]  ( .D(N24), .E(n63), .C(CLK), .RN(n155), .QN(n25) );
  DFEC1 \Addsum_reg[10]  ( .D(N23), .E(n63), .C(CLK), .RN(n155), .QN(n26) );
  DFEC1 \Addsum_reg[9]  ( .D(N22), .E(n63), .C(CLK), .RN(n155), .QN(n27) );
  DFEC1 \Addsum_reg[8]  ( .D(N21), .E(n63), .C(CLK), .RN(n155), .QN(n28) );
  DFEC1 \Addsum_reg[7]  ( .D(N20), .E(n63), .C(CLK), .RN(n155), .QN(n29) );
  DFEC1 \Addsum_reg[6]  ( .D(N19), .E(n63), .C(CLK), .RN(n155), .QN(n30) );
  DFEC1 \Addsum_reg[5]  ( .D(N18), .E(n63), .C(CLK), .RN(n154), .QN(n31) );
  DFEC1 \Addsum_reg[4]  ( .D(N17), .E(n63), .C(CLK), .RN(n155), .QN(n32) );
  DFEC1 \Addsum_reg[3]  ( .D(N16), .E(n63), .C(CLK), .RN(n155), .QN(n33) );
  DFEC1 \Addsum_reg[2]  ( .D(N15), .E(n63), .C(CLK), .RN(n155), .QN(n34) );
  DFEC1 \Addsum_reg[1]  ( .D(N14), .E(n63), .C(CLK), .RN(n155), .QN(n35) );
  DFEC1 \Addsum_reg[0]  ( .D(N13), .E(n63), .C(CLK), .RN(n155), .QN(n36) );
  DFEC1 OUT_STROBE_reg ( .D(n133), .E(n60), .C(CLK), .RN(NRST), .Q(OUT_STROBE)
         );
  INV0 U64 ( .A(n100), .Q(n101) );
  INV0 U65 ( .A(n102), .Q(n103) );
  INV0 U66 ( .A(n104), .Q(n105) );
  INV0 U67 ( .A(n106), .Q(n107) );
  INV0 U68 ( .A(n108), .Q(n109) );
  INV0 U69 ( .A(n110), .Q(n111) );
  INV0 U70 ( .A(n112), .Q(n113) );
  INV0 U71 ( .A(n114), .Q(n115) );
  INV0 U72 ( .A(n116), .Q(n117) );
  INV0 U73 ( .A(n118), .Q(n119) );
  INV0 U74 ( .A(n120), .Q(n121) );
  INV0 U75 ( .A(n122), .Q(n123) );
  INV0 U76 ( .A(n124), .Q(n125) );
  INV0 U77 ( .A(n126), .Q(n127) );
  INV0 U78 ( .A(n128), .Q(n129) );
  CLKIN0 U79 ( .A(n97), .Q(n98) );
  OAI221 U80 ( .A(n61), .B(n18), .C(n36), .D(n62), .Q(n97) );
  INV3 U81 ( .A(n98), .Q(n99) );
  CLKIN0 U82 ( .A(n96), .Q(n100) );
  OAI222 U83 ( .A(n61), .B(n17), .C(n35), .D(n62), .Q(n96) );
  CLKIN0 U84 ( .A(n95), .Q(n102) );
  OAI222 U85 ( .A(n61), .B(n16), .C(n34), .D(n62), .Q(n95) );
  CLKIN0 U86 ( .A(n94), .Q(n104) );
  OAI222 U87 ( .A(n61), .B(n15), .C(n33), .D(n62), .Q(n94) );
  CLKIN0 U88 ( .A(n93), .Q(n106) );
  OAI222 U89 ( .A(n61), .B(n14), .C(n32), .D(n62), .Q(n93) );
  CLKIN0 U90 ( .A(n92), .Q(n108) );
  OAI222 U91 ( .A(n61), .B(n13), .C(n31), .D(n62), .Q(n92) );
  CLKIN0 U92 ( .A(n91), .Q(n110) );
  OAI222 U93 ( .A(n61), .B(n12), .C(n30), .D(n62), .Q(n91) );
  CLKIN0 U94 ( .A(n90), .Q(n112) );
  OAI222 U95 ( .A(n61), .B(n11), .C(n29), .D(n62), .Q(n90) );
  CLKIN0 U96 ( .A(n89), .Q(n114) );
  OAI222 U97 ( .A(n61), .B(n10), .C(n28), .D(n62), .Q(n89) );
  CLKIN0 U98 ( .A(n88), .Q(n116) );
  OAI222 U99 ( .A(n61), .B(n9), .C(n27), .D(n62), .Q(n88) );
  CLKIN0 U100 ( .A(n87), .Q(n118) );
  OAI222 U101 ( .A(n61), .B(n8), .C(n26), .D(n62), .Q(n87) );
  CLKIN0 U102 ( .A(n86), .Q(n120) );
  OAI222 U103 ( .A(n61), .B(n7), .C(n25), .D(n62), .Q(n86) );
  CLKIN0 U104 ( .A(n85), .Q(n122) );
  OAI222 U105 ( .A(n61), .B(n6), .C(n24), .D(n62), .Q(n85) );
  CLKIN0 U106 ( .A(n84), .Q(n124) );
  OAI222 U107 ( .A(n61), .B(n5), .C(n23), .D(n62), .Q(n84) );
  CLKIN0 U108 ( .A(n83), .Q(n126) );
  OAI222 U109 ( .A(n61), .B(n4), .C(n22), .D(n62), .Q(n83) );
  CLKIN0 U110 ( .A(n82), .Q(n128) );
  OAI222 U111 ( .A(n61), .B(n3), .C(n21), .D(n62), .Q(n82) );
  CLKIN0 U112 ( .A(n81), .Q(n130) );
  OAI221 U113 ( .A(n61), .B(n2), .C(n20), .D(n62), .Q(n81) );
  INV3 U114 ( .A(n130), .Q(n131) );
  CLKIN0 U115 ( .A(n19), .Q(n132) );
  INV3 U116 ( .A(n132), .Q(n133) );
  BUF2 U117 ( .A(Add2[0]), .Q(n134) );
  BUF2 U118 ( .A(n80), .Q(n135) );
  NAND20 U119 ( .A(OUT[0]), .B(n157), .Q(n59) );
  BUF2 U120 ( .A(n79), .Q(n136) );
  NAND20 U121 ( .A(OUT[1]), .B(n157), .Q(n58) );
  BUF2 U122 ( .A(n78), .Q(n137) );
  NAND20 U123 ( .A(OUT[2]), .B(n157), .Q(n57) );
  BUF2 U124 ( .A(n77), .Q(n138) );
  NAND20 U125 ( .A(OUT[3]), .B(n157), .Q(n56) );
  BUF2 U126 ( .A(n76), .Q(n139) );
  NAND20 U127 ( .A(OUT[4]), .B(n157), .Q(n55) );
  BUF2 U128 ( .A(n75), .Q(n140) );
  NAND20 U129 ( .A(OUT[5]), .B(n157), .Q(n54) );
  BUF2 U130 ( .A(n74), .Q(n141) );
  NAND20 U131 ( .A(OUT[6]), .B(n157), .Q(n53) );
  BUF2 U132 ( .A(n73), .Q(n142) );
  NAND20 U133 ( .A(OUT[7]), .B(n157), .Q(n52) );
  BUF2 U134 ( .A(n72), .Q(n143) );
  NAND20 U135 ( .A(OUT[8]), .B(n157), .Q(n51) );
  BUF2 U136 ( .A(n71), .Q(n144) );
  NAND20 U137 ( .A(OUT[9]), .B(n157), .Q(n50) );
  BUF2 U138 ( .A(n70), .Q(n145) );
  NAND20 U139 ( .A(OUT[10]), .B(n157), .Q(n49) );
  BUF2 U140 ( .A(n69), .Q(n146) );
  NAND20 U141 ( .A(OUT[11]), .B(n157), .Q(n48) );
  BUF2 U142 ( .A(n68), .Q(n147) );
  NAND20 U143 ( .A(OUT[12]), .B(n157), .Q(n47) );
  BUF2 U144 ( .A(n67), .Q(n148) );
  NAND20 U145 ( .A(OUT[13]), .B(n157), .Q(n46) );
  BUF2 U146 ( .A(n66), .Q(n149) );
  NAND20 U147 ( .A(OUT[14]), .B(n157), .Q(n45) );
  BUF2 U148 ( .A(n65), .Q(n150) );
  NAND20 U149 ( .A(OUT[15]), .B(n157), .Q(n44) );
  BUF2 U150 ( .A(n64), .Q(n151) );
  NAND20 U151 ( .A(OUT[16]), .B(n157), .Q(n43) );
  CLKIN0 U152 ( .A(n40), .Q(n152) );
  INV8 U153 ( .A(n41), .Q(n156) );
  AOI210 U154 ( .A(n40), .B(START), .C(state[1]), .Q(n41) );
  BUF2 U155 ( .A(n42), .Q(n153) );
  INV3 U156 ( .A(n60), .Q(n157) );
  NOR22 U157 ( .A(n40), .B(state[1]), .Q(n63) );
  NAND23 U158 ( .A(state[0]), .B(n153), .Q(n61) );
  NOR21 U159 ( .A(n40), .B(\next_state[1] ), .Q(n60) );
  NAND22 U160 ( .A(n158), .B(n62), .Q(\next_state[1] ) );
  INV3 U161 ( .A(n63), .Q(n158) );
  NAND22 U162 ( .A(n60), .B(n19), .Q(n42) );
  NAND24 U163 ( .A(state[1]), .B(n40), .Q(n62) );
  BUF2 U164 ( .A(NRST), .Q(n154) );
  BUF2 U165 ( .A(NRST), .Q(n155) );
  LOGIC0 U166 ( .Q(n159) );
endmodule


module MatrixMultiplier_DW01_add_0 ( A, B, CI, SUM, CO );
  input [16:0] A;
  input [16:0] B;
  output [16:0] SUM;
  input CI;
  output CO;
  wire   n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n16, n17;
  wire   [16:1] carry;

  XOR30 U1_16 ( .A(A[16]), .B(B[16]), .C(carry[16]), .Q(SUM[16]) );
  ADD31 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(n18)
         );
  ADD31 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(n19)
         );
  ADD31 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(n20)
         );
  ADD31 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(n21)
         );
  ADD31 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(n22)
         );
  ADD31 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(n23)
         );
  ADD31 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(n24) );
  ADD31 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(n25) );
  ADD31 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(n26) );
  ADD31 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(n27) );
  ADD31 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(n28) );
  ADD31 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(n29) );
  ADD31 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(n30) );
  ADD31 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(n31) );
  ADD31 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(n32) );
  XOR20 U1 ( .A(A[0]), .B(B[0]), .Q(SUM[0]) );
  BUF2 U2 ( .A(n32), .Q(SUM[1]) );
  BUF2 U3 ( .A(n31), .Q(SUM[2]) );
  BUF2 U4 ( .A(n30), .Q(SUM[3]) );
  BUF2 U5 ( .A(n29), .Q(SUM[4]) );
  BUF2 U6 ( .A(n28), .Q(SUM[5]) );
  BUF2 U7 ( .A(n27), .Q(SUM[6]) );
  BUF2 U8 ( .A(n26), .Q(SUM[7]) );
  BUF2 U9 ( .A(n25), .Q(SUM[8]) );
  BUF2 U10 ( .A(n24), .Q(SUM[9]) );
  BUF2 U11 ( .A(n23), .Q(SUM[10]) );
  BUF2 U12 ( .A(n22), .Q(SUM[11]) );
  BUF2 U13 ( .A(n21), .Q(SUM[12]) );
  BUF2 U14 ( .A(n20), .Q(SUM[13]) );
  BUF2 U15 ( .A(n19), .Q(SUM[14]) );
  BUF2 U16 ( .A(n18), .Q(SUM[15]) );
  NOR21 U17 ( .A(n16), .B(n17), .Q(carry[1]) );
  INV3 U18 ( .A(B[0]), .Q(n16) );
  INV3 U19 ( .A(A[0]), .Q(n17) );
endmodule


module MatrixMultiplier_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n78, n79, n80, n81, n83, n84,
         n85, n86, n88, n89, n91, n92, n93, n94, n95, n96, n97, n100, n101,
         n102, n103, n104, n105, n107, n108, n109, n110, n111, n112, n113,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283;

  ADD32 U2 ( .A(n218), .B(n15), .CI(n2), .CO(n1), .S(product[14]) );
  ADD32 U3 ( .A(n17), .B(n217), .CI(n3), .CO(n2), .S(product[13]) );
  ADD32 U4 ( .A(n19), .B(n18), .CI(n4), .CO(n3), .S(product[12]) );
  ADD32 U5 ( .A(n20), .B(n23), .CI(n5), .CO(n4), .S(product[11]) );
  ADD32 U6 ( .A(n24), .B(n27), .CI(n6), .CO(n5), .S(product[10]) );
  ADD32 U7 ( .A(n28), .B(n33), .CI(n7), .CO(n6), .S(product[9]) );
  ADD32 U8 ( .A(n34), .B(n40), .CI(n8), .CO(n7), .S(product[8]) );
  ADD32 U9 ( .A(n41), .B(n46), .CI(n9), .CO(n8), .S(product[7]) );
  ADD32 U10 ( .A(n47), .B(n50), .CI(n10), .CO(n9), .S(product[6]) );
  ADD32 U11 ( .A(n51), .B(n53), .CI(n11), .CO(n10), .S(product[5]) );
  ADD32 U12 ( .A(n55), .B(n56), .CI(n12), .CO(n11), .S(product[4]) );
  ADD32 U13 ( .A(n57), .B(n80), .CI(n13), .CO(n12), .S(product[3]) );
  ADD32 U14 ( .A(n105), .B(n112), .CI(n14), .CO(n13), .S(product[2]) );
  ADD22 U15 ( .A(n113), .B(n81), .CO(n14), .S(product[1]) );
  ADD32 U17 ( .A(n83), .B(n21), .CI(n222), .CO(n17), .S(n18) );
  ADD32 U18 ( .A(n221), .B(n84), .CI(n25), .CO(n19), .S(n20) );
  ADD32 U20 ( .A(n29), .B(n226), .CI(n26), .CO(n23), .S(n24) );
  ADD32 U21 ( .A(n91), .B(n31), .CI(n85), .CO(n25), .S(n26) );
  ADD32 U22 ( .A(n35), .B(n216), .CI(n30), .CO(n27), .S(n28) );
  ADD32 U23 ( .A(n86), .B(n92), .CI(n225), .CO(n29), .S(n30) );
  ADD32 U25 ( .A(n39), .B(n42), .CI(n36), .CO(n33), .S(n34) );
  ADD32 U26 ( .A(n229), .B(n93), .CI(n44), .CO(n35), .S(n36) );
  ADD32 U30 ( .A(n45), .B(n48), .CI(n43), .CO(n40), .S(n41) );
  ADD32 U31 ( .A(n88), .B(n100), .CI(n94), .CO(n42), .S(n43) );
  ADD22 U32 ( .A(n78), .B(n107), .CO(n44), .S(n45) );
  ADD32 U33 ( .A(n52), .B(n101), .CI(n49), .CO(n46), .S(n47) );
  ADD32 U34 ( .A(n89), .B(n108), .CI(n95), .CO(n48), .S(n49) );
  ADD32 U35 ( .A(n96), .B(n102), .CI(n54), .CO(n50), .S(n51) );
  ADD22 U36 ( .A(n79), .B(n109), .CO(n52), .S(n53) );
  ADD32 U37 ( .A(n97), .B(n110), .CI(n103), .CO(n54), .S(n55) );
  ADD22 U38 ( .A(n104), .B(n111), .CO(n56), .S(n57) );
  INV1 U166 ( .A(n15), .Q(n217) );
  INV3 U167 ( .A(n1), .Q(product[15]) );
  INV3 U168 ( .A(n265), .Q(n216) );
  INV3 U169 ( .A(n258), .Q(n228) );
  INV3 U170 ( .A(n254), .Q(n218) );
  INV3 U171 ( .A(a[1]), .Q(n230) );
  INV3 U172 ( .A(n260), .Q(n224) );
  INV3 U173 ( .A(n262), .Q(n220) );
  INV3 U174 ( .A(n233), .Q(n226) );
  INV3 U175 ( .A(n277), .Q(n229) );
  INV1 U176 ( .A(n31), .Q(n225) );
  NAND22 U177 ( .A(a[1]), .B(n231), .Q(n256) );
  INV1 U178 ( .A(n21), .Q(n221) );
  INV3 U179 ( .A(n244), .Q(n222) );
  INV3 U180 ( .A(a[3]), .Q(n227) );
  INV3 U181 ( .A(a[5]), .Q(n223) );
  INV3 U182 ( .A(b[0]), .Q(n232) );
  INV3 U183 ( .A(a[7]), .Q(n219) );
  INV3 U184 ( .A(a[0]), .Q(n231) );
  NAND22 U185 ( .A(n224), .B(n268), .Q(n237) );
  NAND22 U186 ( .A(n220), .B(n269), .Q(n247) );
  NAND22 U187 ( .A(n228), .B(n283), .Q(n235) );
  NOR20 U188 ( .A(n231), .B(n232), .Q(product[0]) );
  OAI220 U189 ( .A(n234), .B(n228), .C(n235), .D(n234), .Q(n233) );
  NOR20 U190 ( .A(n224), .B(n232), .Q(n97) );
  OAI220 U191 ( .A(n236), .B(n237), .C(n224), .D(n238), .Q(n96) );
  XNR20 U192 ( .A(n232), .B(n223), .Q(n236) );
  OAI220 U193 ( .A(n238), .B(n237), .C(n224), .D(n239), .Q(n95) );
  XNR20 U194 ( .A(b[1]), .B(a[5]), .Q(n238) );
  OAI220 U195 ( .A(n239), .B(n237), .C(n224), .D(n240), .Q(n94) );
  XNR20 U196 ( .A(b[2]), .B(a[5]), .Q(n239) );
  OAI220 U197 ( .A(n240), .B(n237), .C(n224), .D(n241), .Q(n93) );
  XNR20 U198 ( .A(b[3]), .B(a[5]), .Q(n240) );
  OAI220 U199 ( .A(n241), .B(n237), .C(n224), .D(n242), .Q(n92) );
  XNR20 U200 ( .A(b[4]), .B(a[5]), .Q(n241) );
  OAI220 U201 ( .A(n242), .B(n237), .C(n224), .D(n243), .Q(n91) );
  XNR20 U202 ( .A(b[5]), .B(a[5]), .Q(n242) );
  OAI220 U203 ( .A(n245), .B(n224), .C(n237), .D(n245), .Q(n244) );
  NOR20 U204 ( .A(n220), .B(n232), .Q(n89) );
  OAI220 U205 ( .A(n246), .B(n247), .C(n220), .D(n248), .Q(n88) );
  XNR20 U206 ( .A(n232), .B(n219), .Q(n246) );
  OAI220 U207 ( .A(n249), .B(n247), .C(n220), .D(n250), .Q(n86) );
  OAI220 U208 ( .A(n250), .B(n247), .C(n220), .D(n251), .Q(n85) );
  XNR20 U209 ( .A(b[3]), .B(a[7]), .Q(n250) );
  OAI220 U210 ( .A(n251), .B(n247), .C(n220), .D(n252), .Q(n84) );
  XNR20 U211 ( .A(b[4]), .B(a[7]), .Q(n251) );
  OAI220 U212 ( .A(n252), .B(n247), .C(n220), .D(n253), .Q(n83) );
  XNR20 U213 ( .A(b[5]), .B(a[7]), .Q(n252) );
  OAI220 U214 ( .A(n255), .B(n220), .C(n247), .D(n255), .Q(n254) );
  OAI210 U215 ( .A(b[0]), .B(n230), .C(n256), .Q(n81) );
  OAI210 U216 ( .A(n227), .B(n235), .C(n257), .Q(n80) );
  NAND30 U217 ( .A(n258), .B(n232), .C(a[3]), .Q(n257) );
  OAI210 U218 ( .A(n223), .B(n237), .C(n259), .Q(n79) );
  NAND30 U219 ( .A(n260), .B(n232), .C(a[5]), .Q(n259) );
  OAI210 U220 ( .A(n219), .B(n247), .C(n261), .Q(n78) );
  NAND30 U221 ( .A(n262), .B(n232), .C(a[7]), .Q(n261) );
  XNR20 U222 ( .A(n263), .B(n264), .Q(n39) );
  NOR20 U223 ( .A(n264), .B(n263), .Q(n265) );
  OAI220 U224 ( .A(n248), .B(n247), .C(n220), .D(n249), .Q(n263) );
  XNR20 U225 ( .A(b[2]), .B(a[7]), .Q(n249) );
  XNR20 U226 ( .A(b[1]), .B(a[7]), .Q(n248) );
  OAI220 U227 ( .A(n266), .B(n235), .C(n228), .D(n267), .Q(n264) );
  OAI220 U228 ( .A(n267), .B(n235), .C(n228), .D(n234), .Q(n31) );
  XNR20 U229 ( .A(b[7]), .B(a[3]), .Q(n234) );
  XNR20 U230 ( .A(b[6]), .B(a[3]), .Q(n267) );
  OAI220 U231 ( .A(n243), .B(n237), .C(n224), .D(n245), .Q(n21) );
  XNR20 U232 ( .A(b[7]), .B(a[5]), .Q(n245) );
  XNR20 U233 ( .A(a[4]), .B(n223), .Q(n268) );
  XNR20 U234 ( .A(a[4]), .B(n227), .Q(n260) );
  XNR20 U235 ( .A(b[6]), .B(a[5]), .Q(n243) );
  OAI220 U236 ( .A(n253), .B(n247), .C(n220), .D(n255), .Q(n15) );
  XNR20 U237 ( .A(b[7]), .B(a[7]), .Q(n255) );
  XNR20 U238 ( .A(a[6]), .B(n219), .Q(n269) );
  XNR20 U239 ( .A(a[6]), .B(n223), .Q(n262) );
  XNR20 U240 ( .A(b[6]), .B(a[7]), .Q(n253) );
  OAI220 U241 ( .A(b[0]), .B(n256), .C(n270), .D(n231), .Q(n113) );
  OAI220 U242 ( .A(n270), .B(n256), .C(n271), .D(n231), .Q(n112) );
  XNR20 U243 ( .A(b[1]), .B(a[1]), .Q(n270) );
  OAI220 U244 ( .A(n271), .B(n256), .C(n272), .D(n231), .Q(n111) );
  XNR20 U245 ( .A(b[2]), .B(a[1]), .Q(n271) );
  OAI220 U246 ( .A(n272), .B(n256), .C(n273), .D(n231), .Q(n110) );
  XNR20 U247 ( .A(b[3]), .B(a[1]), .Q(n272) );
  OAI220 U248 ( .A(n273), .B(n256), .C(n274), .D(n231), .Q(n109) );
  XNR20 U249 ( .A(b[4]), .B(a[1]), .Q(n273) );
  OAI220 U250 ( .A(n274), .B(n256), .C(n275), .D(n231), .Q(n108) );
  XNR20 U251 ( .A(b[5]), .B(a[1]), .Q(n274) );
  OAI220 U252 ( .A(n275), .B(n256), .C(n276), .D(n231), .Q(n107) );
  XNR20 U253 ( .A(b[6]), .B(a[1]), .Q(n275) );
  OAI220 U254 ( .A(n231), .B(n276), .C(n256), .D(n276), .Q(n277) );
  XNR20 U255 ( .A(b[7]), .B(a[1]), .Q(n276) );
  NOR20 U256 ( .A(n228), .B(n232), .Q(n105) );
  OAI220 U257 ( .A(n278), .B(n235), .C(n228), .D(n279), .Q(n104) );
  XNR20 U258 ( .A(n232), .B(n227), .Q(n278) );
  OAI220 U259 ( .A(n279), .B(n235), .C(n228), .D(n280), .Q(n103) );
  XNR20 U260 ( .A(b[1]), .B(a[3]), .Q(n279) );
  OAI220 U261 ( .A(n280), .B(n235), .C(n228), .D(n281), .Q(n102) );
  XNR20 U262 ( .A(b[2]), .B(a[3]), .Q(n280) );
  OAI220 U263 ( .A(n281), .B(n235), .C(n228), .D(n282), .Q(n101) );
  XNR20 U264 ( .A(b[3]), .B(a[3]), .Q(n281) );
  OAI220 U265 ( .A(n282), .B(n235), .C(n228), .D(n266), .Q(n100) );
  XNR20 U266 ( .A(b[5]), .B(a[3]), .Q(n266) );
  XNR20 U267 ( .A(a[2]), .B(n227), .Q(n283) );
  XNR20 U268 ( .A(a[2]), .B(n230), .Q(n258) );
  XNR20 U269 ( .A(b[4]), .B(a[3]), .Q(n282) );
endmodule

